// shell for advanced traffic light controller (stretch goal)
// CSE140L   Summer II  2019
// semi-independent operation of east and west straight and left signals
//  see assignment writeup

module traffic_light_controller(
  input clk,
        reset,
        ew_left_sensor,
        ew_str_sensor,		
        ns_sensor,
  output logic[1:0] ew_left_light,     
  		            ew_str_light,	   	
			        ns_light);					  
	

endmodule 